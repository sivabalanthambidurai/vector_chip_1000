//____________________________________________________________________________________________________________________
//file name : lane.sv
//author : sivabalan
//description : This file holds the logic for lane inside the pipeline.
//____________________________________________________________________________________________________________________

module lane (input clk,
             input reset
            );
 
endmodule