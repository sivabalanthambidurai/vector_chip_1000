//____________________________________________________________________________________________________________________
//file name : ifetch_unit.sv
//author : sivabalan
//description : This file holds the logic for instruction fetch unit
//____________________________________________________________________________________________________________________

module ifetch_unit (input clk,
                    input reset
                   ); 
 
endmodule