//____________________________________________________________________________________________________________________
//file name : wb.sv
//author : sivabalan
//description : This file holds the logic for write-back.
//____________________________________________________________________________________________________________________

module wb (input clk,
           input reset
          ); 
 
endmodule