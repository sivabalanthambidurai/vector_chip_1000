//____________________________________________________________________________________________________________________
//file name : crossbar_switch.sv
//author : sivabalan
//description : This file holds the crossbar_switch logic.
//This module is responsible for inter-connecting the different lanes in a core with the core registers
//____________________________________________________________________________________________________________________

module crossbar_switch (input clk,
                        input reset,
                    
                       ); 

endmodule
