//____________________________________________________________________________________________________________________
//file name : stp.sv
//author : sivabalan
//description : This file holds the logic for stp
//____________________________________________________________________________________________________________________

module stp (input clk,
            input reset
           ); 
 
endmodule