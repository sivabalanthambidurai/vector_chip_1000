//____________________________________________________________________________________________________________________
//file name : vector_functional_unit.sv
//author : sivabalan
//description : This file holds the vector functional logic. Vector functional unit holds the following functions
//TODO: 
//____________________________________________________________________________________________________________________

module vector_functional_unit (input clk,
                               input reset

                               );
  
  
endmodule
