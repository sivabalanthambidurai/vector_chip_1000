//____________________________________________________________________________________________________________________
//file name : vector_load_store_unit.sv
//author : sivabalan
//description : This file holds the vector load and store unit. This module is responsible for generating memory read and 
//write request.  
//____________________________________________________________________________________________________________________


module vector_load_store_unit (input clk,
                               input reset

                               );
  
  
endmodule
