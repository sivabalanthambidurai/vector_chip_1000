//____________________________________________________________________________________________________________________
//file name : thread_manager.sv
//author : sivabalan
//description : This file holds the logic for thread manager.
//____________________________________________________________________________________________________________________

module thread_manager (input clk,
                       input reset
                      ); 
 
endmodule