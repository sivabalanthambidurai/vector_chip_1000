//____________________________________________________________________________________________________________________
//file name : core.sv
//author : sivabalan
//description : This file holds the top level core logic.
//____________________________________________________________________________________________________________________

module memory_controller (input clk,
                          input reset,
                    
                          //memory interface
                          input request_t mem_rsp,
                          output request_t mem_req
                       
                          );
  
endmodule
